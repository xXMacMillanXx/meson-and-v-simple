module main

fn main() {
	data := ['one', 'two', 'three', 'four']
	for d in data {
		println('Hello ${d}!')
	}
}
